`default_nettype none

module cpu # (
    parameter BROM_SIZE = 512,
    parameter BROM_INIT = "",

    parameter IMEM_SIZE = 512,
    parameter IMEM_INIT = "",

    parameter DMEM_SIZE = 512,
    parameter DMEM_INIT = "",

    parameter CLK_FREQ = 25000000,
    parameter UART_BAUD = 115200,

    parameter INIT_PC = 32'h10000000,

    parameter USE_BARREL_SHIFTER = 1
) (
    output wire [31:0] o_gpio_out,
    input wire [31:0] i_gpio_in,

`ifdef VERIFICATION
    output wire [31:0] d_regs_out[0:31],
    output wire [31:0] d_finished_instruction,
`endif

    output wire o_tx,
    input wire i_rx,

    input wire i_rst,
    input wire i_clk
);

wire alu_stall;
wire inst_stall;
wire data_stall;
wire stall = alu_stall || inst_stall || data_stall;

wire take_branch;
wire take_jump;
reg [31:0] rd_write;

instruction_t instr_1;
instruction_t instr_2;

wire [31:0] raw_instr;
reg [31:0] pc = INIT_PC - 4;
reg [31:0] next_pc;

wire [31:0] data_addr;
wire [31:0] data_rdata;
wire [31:0] data_wdata;
wire [1:0] data_width;
wire data_we;
wire data_read_en;
wire data_zeroextend;

memory_controller #(
    .BROM_INIT(BROM_INIT),
    .BROM_SIZE(BROM_SIZE),

    .IMEM_INIT(IMEM_INIT),
    .IMEM_SIZE(IMEM_SIZE),

    .DMEM_INIT(DMEM_INIT),
    .DMEM_SIZE(DMEM_SIZE),
    .CLK_FREQ(CLK_FREQ),
    .UART_BAUD(UART_BAUD)
) mem_controller (
    .i_inst_addr(next_pc),
    .o_inst_data(raw_instr),
    .i_inst_re(~stall),
    .o_inst_stall(inst_stall),

    .i_data_addr(data_addr),
    .o_data_data(data_rdata),
    .i_data_data(data_wdata),
    .i_data_width(data_width),
    .i_data_we(data_we),
    .i_data_re(~stall && data_read_en),
    .i_data_zeroextend(data_zeroextend),
    .o_data_stall(data_stall),

    .o_gpio_out(o_gpio_out),
    .i_gpio_in(i_gpio_in),

    .o_tx(o_tx),
    .i_rx(i_rx),

    .i_clk(i_clk),
    .i_rst(i_rst)
);

decode decode (
    .i_instr(raw_instr),
    .i_pc(pc),
    .o_out(instr_1)
);


wire [31:0] rs1_read;
wire [31:0] rs2_read;

// Forwarding
wire fwd1 = ((instr_1.rs1_addr == instr_2.rd_addr) && (instr_2.rd_addr != 0));
wire fwd2 = ((instr_1.rs2_addr == instr_2.rd_addr) && (instr_2.rd_addr != 0));
wire [31:0] rs1 = fwd1 ? rd_write : rs1_read;
wire [31:0] rs2 = fwd2 ? rd_write : rs2_read;

regfile regfile (
    .i_rd_addr(stall ? 0 : instr_2.rd_addr),
    .i_rd_data(rd_write),
    .i_rs1_addr(instr_1.rs1_addr),
    .o_rs1_data(rs1_read),
    .i_rs2_addr(instr_1.rs2_addr),
    .o_rs2_data(rs2_read),

`ifdef VERIFICATION
    .d_regs_out(d_regs_out),
`endif

    .i_clk(i_clk)
);

wire [31:0] alu_A = (instr_1.rs1_pc) ? instr_1.pc : rs1;
wire [31:0] alu_B = (instr_1.rs2_imm) ? instr_1.imm : rs2;

// One cycle delay across ALU
wire [31:0] alu_out;
wire alu_valid;
assign alu_stall = ~alu_valid;
alu #(
    .USE_BARREL_SHIFTER(USE_BARREL_SHIFTER)
) alu (
    .i_op(instr_1.alu_op),
    .i_A(alu_A),
    .i_B(alu_B),
    .o_out(alu_out),
    .i_valid(~stall),
    .o_valid(alu_valid),
    .i_clk(i_clk),
    .i_rst(i_rst)
);

wire branch_out;
assign take_branch = (branch_out && instr_1.branch);
branch_controller branch (
    .i_rs1(rs1),
    .i_rs2(rs2),
    .i_branch_type(instr_1.branch_type),
    .o_take_branch(branch_out)
);

assign take_jump = instr_1.jump;

assign data_wdata = rs2;
assign data_addr = (rs1 + instr_1.imm);
assign data_width = instr_1.loadstore[1:0];
assign data_we = ~stall && (instr_1.loadstore > 4);
assign data_read_en = ~stall && ((instr_1.loadstore > 0) && (instr_1.loadstore < 4));
assign data_zeroextend = instr_1.load_zeroextend;

always_comb begin
    if (instr_2.jump) begin
        rd_write = instr_2.pc + 4;
    end
    else if ((instr_2.loadstore > 0) && (instr_2.loadstore < 4)) begin
        rd_write = data_rdata;
    end
    else begin
        rd_write = alu_out;
    end
end

always_comb begin
    if (i_rst) begin
        next_pc = INIT_PC;
    end
    else if (stall) begin
        next_pc = pc;
    end
    else if (take_jump | take_branch) begin
        next_pc = alu_A + alu_B;
    end
    else begin
        next_pc = pc + 4;
    end
end

initial begin
    instr_1 = 0;
    instr_2 = 0;
end

always_ff @(posedge i_clk) begin
    if (~stall) begin
        instr_2 <= i_rst ? 0 : instr_1;
        pc <= next_pc;
    end
end

`ifdef VERIFICATION
    assign d_finished_instruction = instr_2.inst_raw[32] == 1 ? (instr_2.inst_raw[31:0]) : 0;
`endif

endmodule
