`default_nettype none

module top (
    input wire i_clk
);

endmodule
